package exn_pkg;
endpackage